// Module for Instruction Memory

module memory(prog_counter, instruction);

	reg [31:0] REGISTER[0:7];									// 8 32-bit memory register

	input [2:0] prog_counter; 									// 3 bit program counter as input
	output wire [31:0] instruction;								// 32 bit instruction as output

	initial
		begin
			REGISTER[0] = 32'b00100000000001000011010001010110;	// 001000 00000 00100  (0011 0100 0101 0110)
			REGISTER[1] = 32'b00100000000001011111111111111111;	// 001000 00000 00101  (1111 1111 1111 1111)
			REGISTER[2] = 32'b00000000101001000011000000010000;	// 000000 00101 00100 00110 00000 010000 
			REGISTER[3] = 32'b00100000000000110000000000000111;	// 001000 00000 00011  (0000 0000 0000 0111)
			REGISTER[4] = 32'b00000000110000110011000000000100;	// 000000 00110 00011 00110 00000 000100
			REGISTER[5] = 32'b00000000000000110001100001000010; // 000000 00000 00011 00011 00001 000010
			REGISTER[6] = 32'b10001100100001011001101010111100; // 100011 00100 00101 (1001 1010 1011 1100)
			REGISTER[7] = 32'b00001000000100100011010001010110; // 000010 (00 0001 0010 0011 0100 0101 0110)
		end

	assign instruction = REGISTER[prog_counter];				// Multiplexer to choose the instruction from the program counter

endmodule